
// Alguma coisa pra teste...

module ok(a , b, c);

input a;// sinal de entrada
input b;
output c;

wire tmp, af, gr;

not #2(tmp, a);

and(c, tmp, af ,);

endmodule



