
// Alguma coisa pra teste

module ok(a , b, c);

input a;// sinal de entrada

input b;

output c;

and(a, x, y);

endmodule