
/*

blah blah
blah

*/

module multiline();

/*nada*/

  /* mais nada */

/**/

  wire w;

/*  */

/*//*/

/*/////*/

/* // */

/* ///// */

/*  //
    //
        */

endmodule /* final */

