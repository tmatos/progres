
// Alguma coisa pra teste

module ok(a , b, c);

input a;// sinal de entrada
input b;
output c;

wire tmp;

not(tmp, a); and(a, x, y);

endmodule