
// Alguma coisa pra teste, (bugada)

module ok(a , ok, c);

input a;// sinal de entrada

and(a, x, y);

endmodule