
// Alguma coisa pra teste

module ok(a , b, c);

input a;// sinal de entrada
input b;
output c;

wire tmp;

not(c, a); and(a, x, y);

endmodule