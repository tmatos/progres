
// Alguma coisa pra teste

module ok(a, b, c)

in a;// sinal de entrada

and(a, x, y);

end module