
// Alguma coisa pra teste

module ok(a , b, c);

input a;// sinal de entrada

and(a, x, y);

endmodule