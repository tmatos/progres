
module top();

endmodule
